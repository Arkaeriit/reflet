/*
 * This rom is made from the proram test_instruction.asm.
 * It is meant to test most instructions.
 */
module rom8(input clk, input enable, input [14-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            9'h0 : data_reg <= 16'h5341;
            9'h1 : data_reg <= 16'h4D52;
            9'h2 : data_reg <= 16'h2D3C;
            9'h3 : data_reg <= 16'h2C3B;
            9'h4 : data_reg <= 16'h3D10;
            9'h5 : data_reg <= 16'h3C12;
            9'h6 : data_reg <= 16'h0000;
            9'h7 : data_reg <= 16'h0000;
            9'h8 : data_reg <= 16'h4C12;
            9'h9 : data_reg <= 16'h3E4E;
            9'hA : data_reg <= 16'h039C;
            9'hB : data_reg <= 16'h4C13;
            9'hC : data_reg <= 16'h4E08;
            9'hD : data_reg <= 16'h3CF0;
            9'hE : data_reg <= 16'h3D2B;
            9'hF : data_reg <= 16'h3F2C;
            9'h10 : data_reg <= 16'h2D3C;
            9'h11 : data_reg <= 16'h2C3B;
            9'h12 : data_reg <= 16'h3D10;
            9'h13 : data_reg <= 16'h3C12;
            9'h14 : data_reg <= 16'h0000;
            9'h15 : data_reg <= 16'h0000;
            9'h16 : data_reg <= 16'h4C12;
            9'h17 : data_reg <= 16'h3E4E;
            9'h18 : data_reg <= 16'h0328;
            9'h19 : data_reg <= 16'h4C13;
            9'h1A : data_reg <= 16'h4E08;
            9'h1B : data_reg <= 16'h3CF0;
            9'h1C : data_reg <= 16'h3D2B;
            9'h1D : data_reg <= 16'h3E2C;
            9'h1E : data_reg <= 16'h9000;
            9'h1F : data_reg <= 16'h0014;
            9'h20 : data_reg <= 16'h8000;
            9'h21 : data_reg <= 16'hE921;
            9'h22 : data_reg <= 16'h4912;
            9'h23 : data_reg <= 16'h0D39;
            9'h24 : data_reg <= 16'h2D3C;
            9'h25 : data_reg <= 16'h2C3B;
            9'h26 : data_reg <= 16'h3D10;
            9'h27 : data_reg <= 16'h3C12;
            9'h28 : data_reg <= 16'h0000;
            9'h29 : data_reg <= 16'h0000;
            9'h2A : data_reg <= 16'h4C12;
            9'h2B : data_reg <= 16'h3E4E;
            9'h2C : data_reg <= 16'h003C;
            9'h2D : data_reg <= 16'h4C13;
            9'h2E : data_reg <= 16'h4E08;
            9'h2F : data_reg <= 16'h3CF0;
            9'h30 : data_reg <= 16'h3D2B;
            9'h31 : data_reg <= 16'hF02C;
            9'h32 : data_reg <= 16'h3C31;
            9'h33 : data_reg <= 16'h3B2D;
            9'h34 : data_reg <= 16'h102C;
            9'h35 : data_reg <= 16'h123D;
            9'h36 : data_reg <= 16'h003C;
            9'h37 : data_reg <= 16'h0000;
            9'h38 : data_reg <= 16'h0000;
            9'h39 : data_reg <= 16'h4C12;
            9'h3A : data_reg <= 16'h3E4E;
            9'h3B : data_reg <= 16'h003E;
            9'h3C : data_reg <= 16'h4C13;
            9'h3D : data_reg <= 16'h4E08;
            9'h3E : data_reg <= 16'h3CF0;
            9'h3F : data_reg <= 16'h3D2B;
            9'h40 : data_reg <= 16'hF02C;
            9'h41 : data_reg <= 16'h1032;
            9'h42 : data_reg <= 16'h1033;
            9'h43 : data_reg <= 16'h12E1;
            9'h44 : data_reg <= 16'h3141;
            9'h45 : data_reg <= 16'h4311;
            9'h46 : data_reg <= 16'h2233;
            9'h47 : data_reg <= 16'h01C3;
            9'h48 : data_reg <= 16'h2D3C;
            9'h49 : data_reg <= 16'h2C3B;
            9'h4A : data_reg <= 16'h3D10;
            9'h4B : data_reg <= 16'h3C12;
            9'h4C : data_reg <= 16'h0000;
            9'h4D : data_reg <= 16'h0000;
            9'h4E : data_reg <= 16'h4C12;
            9'h4F : data_reg <= 16'h3E4E;
            9'h50 : data_reg <= 16'h0085;
            9'h51 : data_reg <= 16'h4C13;
            9'h52 : data_reg <= 16'h4E08;
            9'h53 : data_reg <= 16'h3CF0;
            9'h54 : data_reg <= 16'h3D2B;
            9'h55 : data_reg <= 16'h092C;
            9'h56 : data_reg <= 16'h3C0D;
            9'h57 : data_reg <= 16'h3B2D;
            9'h58 : data_reg <= 16'h102C;
            9'h59 : data_reg <= 16'h123D;
            9'h5A : data_reg <= 16'h003C;
            9'h5B : data_reg <= 16'h0000;
            9'h5C : data_reg <= 16'h0000;
            9'h5D : data_reg <= 16'h4C12;
            9'h5E : data_reg <= 16'h3E4E;
            9'h5F : data_reg <= 16'h003C;
            9'h60 : data_reg <= 16'h4C13;
            9'h61 : data_reg <= 16'h4E08;
            9'h62 : data_reg <= 16'h3CF0;
            9'h63 : data_reg <= 16'h3D2B;
            9'h64 : data_reg <= 16'hF02C;
            9'h65 : data_reg <= 16'h3C31;
            9'h66 : data_reg <= 16'h3B2D;
            9'h67 : data_reg <= 16'h102C;
            9'h68 : data_reg <= 16'h123D;
            9'h69 : data_reg <= 16'h003C;
            9'h6A : data_reg <= 16'h0000;
            9'h6B : data_reg <= 16'h0000;
            9'h6C : data_reg <= 16'h4C12;
            9'h6D : data_reg <= 16'h3E4E;
            9'h6E : data_reg <= 16'h003E;
            9'h6F : data_reg <= 16'h4C13;
            9'h70 : data_reg <= 16'h4E08;
            9'h71 : data_reg <= 16'h3CF0;
            9'h72 : data_reg <= 16'h3D2B;
            9'h73 : data_reg <= 16'hF02C;
            9'h74 : data_reg <= 16'h1032;
            9'h75 : data_reg <= 16'hF133;
            9'h76 : data_reg <= 16'h120F;
            9'h77 : data_reg <= 16'h3141;
            9'h78 : data_reg <= 16'h4311;
            9'h79 : data_reg <= 16'h2233;
            9'h7A : data_reg <= 16'h01C3;
            9'h7B : data_reg <= 16'h2D3C;
            9'h7C : data_reg <= 16'h2C3B;
            9'h7D : data_reg <= 16'h3D10;
            9'h7E : data_reg <= 16'h3C12;
            9'h7F : data_reg <= 16'h0000;
            9'h80 : data_reg <= 16'h0000;
            9'h81 : data_reg <= 16'h4C12;
            9'h82 : data_reg <= 16'h3E4E;
            9'h83 : data_reg <= 16'h00EB;
            9'h84 : data_reg <= 16'h4C13;
            9'h85 : data_reg <= 16'h4E08;
            9'h86 : data_reg <= 16'h3CF0;
            9'h87 : data_reg <= 16'h3D2B;
            9'h88 : data_reg <= 16'h092C;
            9'h89 : data_reg <= 16'h3C0D;
            9'h8A : data_reg <= 16'h3B2D;
            9'h8B : data_reg <= 16'h102C;
            9'h8C : data_reg <= 16'h123D;
            9'h8D : data_reg <= 16'h003C;
            9'h8E : data_reg <= 16'h0000;
            9'h8F : data_reg <= 16'h0000;
            9'h90 : data_reg <= 16'h4C12;
            9'h91 : data_reg <= 16'h3E4E;
            9'h92 : data_reg <= 16'h003C;
            9'h93 : data_reg <= 16'h4C13;
            9'h94 : data_reg <= 16'h4E08;
            9'h95 : data_reg <= 16'h3CF0;
            9'h96 : data_reg <= 16'h3D2B;
            9'h97 : data_reg <= 16'hF02C;
            9'h98 : data_reg <= 16'h3C39;
            9'h99 : data_reg <= 16'h3B2D;
            9'h9A : data_reg <= 16'h102C;
            9'h9B : data_reg <= 16'h123D;
            9'h9C : data_reg <= 16'h003C;
            9'h9D : data_reg <= 16'h0000;
            9'h9E : data_reg <= 16'h0000;
            9'h9F : data_reg <= 16'h4C12;
            9'hA0 : data_reg <= 16'h3E4E;
            9'hA1 : data_reg <= 16'h0042;
            9'hA2 : data_reg <= 16'h4C13;
            9'hA3 : data_reg <= 16'h4E08;
            9'hA4 : data_reg <= 16'h3CF0;
            9'hA5 : data_reg <= 16'h3D2B;
            9'hA6 : data_reg <= 16'h3A2C;
            9'hA7 : data_reg <= 16'h3116;
            9'hA8 : data_reg <= 16'h0C2A;
            9'hA9 : data_reg <= 16'h2D3C;
            9'hAA : data_reg <= 16'h2C3B;
            9'hAB : data_reg <= 16'h3D10;
            9'hAC : data_reg <= 16'h3C12;
            9'hAD : data_reg <= 16'h0000;
            9'hAE : data_reg <= 16'h0000;
            9'hAF : data_reg <= 16'h4C12;
            9'hB0 : data_reg <= 16'h3E4E;
            9'hB1 : data_reg <= 16'h0C80;
            9'hB2 : data_reg <= 16'h4C13;
            9'hB3 : data_reg <= 16'h4E08;
            9'hB4 : data_reg <= 16'h3CF0;
            9'hB5 : data_reg <= 16'h3D2B;
            9'hB6 : data_reg <= 16'h322C;
            9'hB7 : data_reg <= 16'h3122;
            9'hB8 : data_reg <= 16'h0C2A;
            9'hB9 : data_reg <= 16'h3C14;
            9'hBA : data_reg <= 16'hAC10;
            9'hBB : data_reg <= 16'h1A3C;
            9'hBC : data_reg <= 16'h317C;
            9'hBD : data_reg <= 16'h3C14;
            9'hBE : data_reg <= 16'hAC10;
            9'hBF : data_reg <= 16'h1F3C;
            9'hC0 : data_reg <= 16'h417C;
            9'hC1 : data_reg <= 16'h2A31;
            9'hC2 : data_reg <= 16'h140C;
            9'hC3 : data_reg <= 16'h163C;
            9'hC4 : data_reg <= 16'h3CAC;
            9'hC5 : data_reg <= 16'h7C14;
            9'hC6 : data_reg <= 16'h1432;
            9'hC7 : data_reg <= 16'h1C3C;
            9'hC8 : data_reg <= 16'h3CAC;
            9'hC9 : data_reg <= 16'h7C18;
            9'hCA : data_reg <= 16'h3152;
            9'hCB : data_reg <= 16'h0C2A;
            9'hCC : data_reg <= 16'h3C14;
            9'hCD : data_reg <= 16'hAC13;
            9'hCE : data_reg <= 16'h123C;
            9'hCF : data_reg <= 16'h527C;
            9'hD0 : data_reg <= 16'h2A31;
            9'hD1 : data_reg <= 16'h140C;
            9'hD2 : data_reg <= 16'h1A3C;
            9'hD3 : data_reg <= 16'h3CAC;
            9'hD4 : data_reg <= 16'h7C1A;
            9'hD5 : data_reg <= 16'h1432;
            9'hD6 : data_reg <= 16'h153C;
            9'hD7 : data_reg <= 16'h3CAC;
            9'hD8 : data_reg <= 16'h7C15;
            9'hD9 : data_reg <= 16'h3162;
            9'hDA : data_reg <= 16'h0C2A;
            9'hDB : data_reg <= 16'h6212;
            9'hDC : data_reg <= 16'h2A31;
            9'hDD : data_reg <= 16'h140C;
            9'hDE : data_reg <= 16'h1A3C;
            9'hDF : data_reg <= 16'h3CAC;
            9'hE0 : data_reg <= 16'h7C1A;
            9'hE1 : data_reg <= 16'h1432;
            9'hE2 : data_reg <= 16'h153C;
            9'hE3 : data_reg <= 16'h3CAC;
            9'hE4 : data_reg <= 16'h7C15;
            9'hE5 : data_reg <= 16'h3172;
            9'hE6 : data_reg <= 16'h0C2A;
            9'hE7 : data_reg <= 16'h331D;
            9'hE8 : data_reg <= 16'h831E;
            9'hE9 : data_reg <= 16'h2A31;
            9'hEA : data_reg <= 16'h920C;
            9'hEB : data_reg <= 16'h2A31;
            9'hEC : data_reg <= 16'h110C;
            9'hED : data_reg <= 16'h1732;
            9'hEE : data_reg <= 16'h31A2;
            9'hEF : data_reg <= 16'h0C2A;
            9'hF0 : data_reg <= 16'hB216;
            9'hF1 : data_reg <= 16'h2A31;
            9'hF2 : data_reg <= 16'h110C;
            9'hF3 : data_reg <= 16'h1131;
            9'hF4 : data_reg <= 16'h3CC1;
            9'hF5 : data_reg <= 16'h3B2D;
            9'hF6 : data_reg <= 16'h102C;
            9'hF7 : data_reg <= 16'h123D;
            9'hF8 : data_reg <= 16'h003C;
            9'hF9 : data_reg <= 16'h0000;
            9'hFA : data_reg <= 16'h0000;
            9'hFB : data_reg <= 16'h4C12;
            9'hFC : data_reg <= 16'h3E4E;
            9'hFD : data_reg <= 16'h0222;
            9'hFE : data_reg <= 16'h4C13;
            9'hFF : data_reg <= 16'h4E08;
            9'h100 : data_reg <= 16'h3CF0;
            9'h101 : data_reg <= 16'h3D2B;
            9'h102 : data_reg <= 16'h092C;
            9'h103 : data_reg <= 16'h2D3C;
            9'h104 : data_reg <= 16'h2C3B;
            9'h105 : data_reg <= 16'h3D10;
            9'h106 : data_reg <= 16'h3C12;
            9'h107 : data_reg <= 16'h0000;
            9'h108 : data_reg <= 16'h0000;
            9'h109 : data_reg <= 16'h4C12;
            9'h10A : data_reg <= 16'h3E4E;
            9'h10B : data_reg <= 16'h0322;
            9'h10C : data_reg <= 16'h4C13;
            9'h10D : data_reg <= 16'h4E08;
            9'h10E : data_reg <= 16'h3CF0;
            9'h10F : data_reg <= 16'h3D2B;
            9'h110 : data_reg <= 16'h3E2C;
            9'h111 : data_reg <= 16'hC110;
            9'h112 : data_reg <= 16'h2D3C;
            9'h113 : data_reg <= 16'h2C3B;
            9'h114 : data_reg <= 16'h3D10;
            9'h115 : data_reg <= 16'h3C12;
            9'h116 : data_reg <= 16'h0000;
            9'h117 : data_reg <= 16'h0000;
            9'h118 : data_reg <= 16'h4C12;
            9'h119 : data_reg <= 16'h3E4E;
            9'h11A : data_reg <= 16'h0322;
            9'h11B : data_reg <= 16'h4C13;
            9'h11C : data_reg <= 16'h4E08;
            9'h11D : data_reg <= 16'h3CF0;
            9'h11E : data_reg <= 16'h3D2B;
            9'h11F : data_reg <= 16'h092C;
            9'h120 : data_reg <= 16'hD111;
            9'h121 : data_reg <= 16'h2D3C;
            9'h122 : data_reg <= 16'h2C3B;
            9'h123 : data_reg <= 16'h3D10;
            9'h124 : data_reg <= 16'h3C12;
            9'h125 : data_reg <= 16'h0000;
            9'h126 : data_reg <= 16'h0000;
            9'h127 : data_reg <= 16'h4C12;
            9'h128 : data_reg <= 16'h3E4E;
            9'h129 : data_reg <= 16'h0322;
            9'h12A : data_reg <= 16'h4C13;
            9'h12B : data_reg <= 16'h4E08;
            9'h12C : data_reg <= 16'h3CF0;
            9'h12D : data_reg <= 16'h3D2B;
            9'h12E : data_reg <= 16'h092C;
            9'h12F : data_reg <= 16'hD110;
            9'h130 : data_reg <= 16'h2D3C;
            9'h131 : data_reg <= 16'h2C3B;
            9'h132 : data_reg <= 16'h3D10;
            9'h133 : data_reg <= 16'h3C12;
            9'h134 : data_reg <= 16'h0000;
            9'h135 : data_reg <= 16'h0000;
            9'h136 : data_reg <= 16'h4C12;
            9'h137 : data_reg <= 16'h3E4E;
            9'h138 : data_reg <= 16'h0298;
            9'h139 : data_reg <= 16'h4C13;
            9'h13A : data_reg <= 16'h4E08;
            9'h13B : data_reg <= 16'h3CF0;
            9'h13C : data_reg <= 16'h3D2B;
            9'h13D : data_reg <= 16'h092C;
            9'h13E : data_reg <= 16'h2D3C;
            9'h13F : data_reg <= 16'h2C3B;
            9'h140 : data_reg <= 16'h3D10;
            9'h141 : data_reg <= 16'h3C12;
            9'h142 : data_reg <= 16'h0000;
            9'h143 : data_reg <= 16'h0000;
            9'h144 : data_reg <= 16'h4C12;
            9'h145 : data_reg <= 16'h3E4E;
            9'h146 : data_reg <= 16'h0322;
            9'h147 : data_reg <= 16'h4C13;
            9'h148 : data_reg <= 16'h4E08;
            9'h149 : data_reg <= 16'h3CF0;
            9'h14A : data_reg <= 16'h3D2B;
            9'h14B : data_reg <= 16'h3E2C;
            9'h14C : data_reg <= 16'h3C14;
            9'h14D : data_reg <= 16'hAC15;
            9'h14E : data_reg <= 16'h1A3C;
            9'h14F : data_reg <= 16'hEF7C;
            9'h150 : data_reg <= 16'hFF10;
            9'h151 : data_reg <= 16'h2A31;
            9'h152 : data_reg <= 16'h140C;
            9'h153 : data_reg <= 16'h153C;
            9'h154 : data_reg <= 16'h3CAC;
            9'h155 : data_reg <= 16'h7C10;
            9'h156 : data_reg <= 16'h100B;
            9'h157 : data_reg <= 16'h310A;
            9'h158 : data_reg <= 16'h0C2A;
            9'h159 : data_reg <= 16'h3C14;
            9'h15A : data_reg <= 16'hAC10;
            9'h15B : data_reg <= 16'h1D3C;
            9'h15C : data_reg <= 16'h087C;
            9'h15D : data_reg <= 16'h2A31;
            9'h15E : data_reg <= 16'h3C0C;
            9'h15F : data_reg <= 16'h3B2D;
            9'h160 : data_reg <= 16'h102C;
            9'h161 : data_reg <= 16'h123D;
            9'h162 : data_reg <= 16'h003C;
            9'h163 : data_reg <= 16'h0000;
            9'h164 : data_reg <= 16'h0000;
            9'h165 : data_reg <= 16'h4C12;
            9'h166 : data_reg <= 16'h3E4E;
            9'h167 : data_reg <= 16'h0323;
            9'h168 : data_reg <= 16'h4C13;
            9'h169 : data_reg <= 16'h4E08;
            9'h16A : data_reg <= 16'h3CF0;
            9'h16B : data_reg <= 16'h3D2B;
            9'h16C : data_reg <= 16'h0C2C;
            9'h16D : data_reg <= 16'h3111;
            9'h16E : data_reg <= 16'hC111;
            9'h16F : data_reg <= 16'h2D3C;
            9'h170 : data_reg <= 16'h2C3B;
            9'h171 : data_reg <= 16'h3D10;
            9'h172 : data_reg <= 16'h3C12;
            9'h173 : data_reg <= 16'h0000;
            9'h174 : data_reg <= 16'h0000;
            9'h175 : data_reg <= 16'h4C12;
            9'h176 : data_reg <= 16'h3E4E;
            9'h177 : data_reg <= 16'h0322;
            9'h178 : data_reg <= 16'h4C13;
            9'h179 : data_reg <= 16'h4E08;
            9'h17A : data_reg <= 16'h3CF0;
            9'h17B : data_reg <= 16'h3D2B;
            9'h17C : data_reg <= 16'h012C;
            9'h17D : data_reg <= 16'h1809;
            9'h17E : data_reg <= 16'h314F;
            9'h17F : data_reg <= 16'h2D3C;
            9'h180 : data_reg <= 16'h2C3B;
            9'h181 : data_reg <= 16'h3D10;
            9'h182 : data_reg <= 16'h3C12;
            9'h183 : data_reg <= 16'h0000;
            9'h184 : data_reg <= 16'h0000;
            9'h185 : data_reg <= 16'h4C12;
            9'h186 : data_reg <= 16'h3E4E;
            9'h187 : data_reg <= 16'hFFFF;
            9'h188 : data_reg <= 16'h4C13;
            9'h189 : data_reg <= 16'h4E08;
            9'h18A : data_reg <= 16'h3CF0;
            9'h18B : data_reg <= 16'h3D2B;
            9'h18C : data_reg <= 16'h032C;
            9'h18D : data_reg <= 16'h10E1;
            9'h18E : data_reg <= 16'h03F1;
            9'h18F : data_reg <= 16'h2A31;
            9'h190 : data_reg <= 16'h0D0C;
            9'h191 : data_reg <= 16'h1A0E;
            9'h192 : data_reg <= 16'h2A31;
            9'h193 : data_reg <= 16'h0D0C;
            9'h194 : data_reg <= 16'h2D3C;
            9'h195 : data_reg <= 16'h2C3B;
            9'h196 : data_reg <= 16'h3D10;
            9'h197 : data_reg <= 16'h3C12;
            9'h198 : data_reg <= 16'h0000;
            9'h199 : data_reg <= 16'h0000;
            9'h19A : data_reg <= 16'h4C12;
            9'h19B : data_reg <= 16'h3E4E;
            9'h19C : data_reg <= 16'h0040;
            9'h19D : data_reg <= 16'h4C13;
            9'h19E : data_reg <= 16'h4E08;
            9'h19F : data_reg <= 16'h3CF0;
            9'h1A0 : data_reg <= 16'h3D2B;
            9'h1A1 : data_reg <= 16'hF02C;
            9'h1A2 : data_reg <= 16'h3C3F;
            9'h1A3 : data_reg <= 16'h3B2D;
            9'h1A4 : data_reg <= 16'h102C;
            9'h1A5 : data_reg <= 16'h123D;
            9'h1A6 : data_reg <= 16'h003C;
            9'h1A7 : data_reg <= 16'h0000;
            9'h1A8 : data_reg <= 16'h0000;
            9'h1A9 : data_reg <= 16'h4C12;
            9'h1AA : data_reg <= 16'h3E4E;
            9'h1AB : data_reg <= 16'h0048;
            9'h1AC : data_reg <= 16'h4C13;
            9'h1AD : data_reg <= 16'h4E08;
            9'h1AE : data_reg <= 16'h3CF0;
            9'h1AF : data_reg <= 16'h3D2B;
            9'h1B0 : data_reg <= 16'h0C2C;
            9'h1B1 : data_reg <= 16'h2D3C;
            9'h1B2 : data_reg <= 16'h2C3B;
            9'h1B3 : data_reg <= 16'h3D10;
            9'h1B4 : data_reg <= 16'h3C12;
            9'h1B5 : data_reg <= 16'h0000;
            9'h1B6 : data_reg <= 16'h0000;
            9'h1B7 : data_reg <= 16'h4C12;
            9'h1B8 : data_reg <= 16'h3E4E;
            9'h1B9 : data_reg <= 16'h0113;
            9'h1BA : data_reg <= 16'h4C13;
            9'h1BB : data_reg <= 16'h4E08;
            9'h1BC : data_reg <= 16'h3CF0;
            9'h1BD : data_reg <= 16'h3D2B;
            9'h1BE : data_reg <= 16'h0C2C;
            9'h1BF : data_reg <= 16'h2D3C;
            9'h1C0 : data_reg <= 16'h2C3B;
            9'h1C1 : data_reg <= 16'h3D10;
            9'h1C2 : data_reg <= 16'h3C12;
            9'h1C3 : data_reg <= 16'h0000;
            9'h1C4 : data_reg <= 16'h0000;
            9'h1C5 : data_reg <= 16'h4C12;
            9'h1C6 : data_reg <= 16'h3E4E;
            9'h1C7 : data_reg <= 16'h00AD;
            9'h1C8 : data_reg <= 16'h4C13;
            9'h1C9 : data_reg <= 16'h4E08;
            9'h1CA : data_reg <= 16'h3CF0;
            9'h1CB : data_reg <= 16'h3D2B;
            9'h1CC : data_reg <= 16'h0C2C;
            9'h1CD : data_reg <= 16'h000E;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
