module rom04(input clk, input enable, input [14-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            14'h0 : data_reg <= 16'h5341;
            14'h1 : data_reg <= 16'h4D52;
            14'h2 : data_reg <= 16'h1C28;
            14'h3 : data_reg <= 16'h9C0D;
            14'h4 : data_reg <= 16'h6D8C;
            14'h5 : data_reg <= 16'h221D;
            14'h6 : data_reg <= 16'h5D8C;
            14'h7 : data_reg <= 16'h1C1D;
            14'h8 : data_reg <= 16'h1B0D;
            14'h9 : data_reg <= 16'h280C;
            14'hA : data_reg <= 16'h0D1C;
            14'hB : data_reg <= 16'h8C9C;
            14'hC : data_reg <= 16'h1D6D;
            14'hD : data_reg <= 16'h8C22;
            14'hE : data_reg <= 16'h1D5D;
            14'hF : data_reg <= 16'h221D;
            14'h10 : data_reg <= 16'h001C;
            14'h11 : data_reg <= 16'h3C22;
            14'h12 : data_reg <= 16'h1E3E;
            14'h13 : data_reg <= 16'h044A;
            14'h14 : data_reg <= 16'h3C23;
            14'h15 : data_reg <= 16'h3EE5;
            14'h16 : data_reg <= 16'h1CD0;
            14'h17 : data_reg <= 16'h1D0B;
            14'h18 : data_reg <= 16'h1F0C;
            14'h19 : data_reg <= 16'h0D1C;
            14'h1A : data_reg <= 16'h0C1B;
            14'h1B : data_reg <= 16'h1C28;
            14'h1C : data_reg <= 16'h9C0D;
            14'h1D : data_reg <= 16'h6D8C;
            14'h1E : data_reg <= 16'h221D;
            14'h1F : data_reg <= 16'h5D8C;
            14'h20 : data_reg <= 16'h1D1D;
            14'h21 : data_reg <= 16'h1C22;
            14'h22 : data_reg <= 16'h3C22;
            14'h23 : data_reg <= 16'h1E3E;
            14'h24 : data_reg <= 16'h03BE;
            14'h25 : data_reg <= 16'h3C23;
            14'h26 : data_reg <= 16'h3EE5;
            14'h27 : data_reg <= 16'h1CD0;
            14'h28 : data_reg <= 16'h1D0B;
            14'h29 : data_reg <= 16'h1E0C;
            14'h2A : data_reg <= 16'h9000;
            14'h2B : data_reg <= 16'h0014;
            14'h2C : data_reg <= 16'h8000;
            14'h2D : data_reg <= 16'hC901;
            14'h2E : data_reg <= 16'h221C;
            14'h2F : data_reg <= 16'h1939;
            14'h30 : data_reg <= 16'hE20C;
            14'h31 : data_reg <= 16'h0D1C;
            14'h32 : data_reg <= 16'h0C1B;
            14'h33 : data_reg <= 16'h1C28;
            14'h34 : data_reg <= 16'h9C0D;
            14'h35 : data_reg <= 16'h6D8C;
            14'h36 : data_reg <= 16'h221D;
            14'h37 : data_reg <= 16'h5D8C;
            14'h38 : data_reg <= 16'h1D1D;
            14'h39 : data_reg <= 16'h1C22;
            14'h3A : data_reg <= 16'h3C22;
            14'h3B : data_reg <= 16'h1E3E;
            14'h3C : data_reg <= 16'h0054;
            14'h3D : data_reg <= 16'h3C23;
            14'h3E : data_reg <= 16'h3EE5;
            14'h3F : data_reg <= 16'h1CD0;
            14'h40 : data_reg <= 16'h1D0B;
            14'h41 : data_reg <= 16'hD00C;
            14'h42 : data_reg <= 16'h1C11;
            14'h43 : data_reg <= 16'h1B0D;
            14'h44 : data_reg <= 16'h280C;
            14'h45 : data_reg <= 16'h0D1C;
            14'h46 : data_reg <= 16'h8C9C;
            14'h47 : data_reg <= 16'h1D6D;
            14'h48 : data_reg <= 16'h8C22;
            14'h49 : data_reg <= 16'h1D5D;
            14'h4A : data_reg <= 16'h221D;
            14'h4B : data_reg <= 16'h001C;
            14'h4C : data_reg <= 16'h3C22;
            14'h4D : data_reg <= 16'h1E3E;
            14'h4E : data_reg <= 16'h0056;
            14'h4F : data_reg <= 16'h3C23;
            14'h50 : data_reg <= 16'h3EE5;
            14'h51 : data_reg <= 16'h1CD0;
            14'h52 : data_reg <= 16'h1D0B;
            14'h53 : data_reg <= 16'hD00C;
            14'h54 : data_reg <= 16'h2012;
            14'h55 : data_reg <= 16'h2013;
            14'h56 : data_reg <= 16'h1CC1;
            14'h57 : data_reg <= 16'h3122;
            14'h58 : data_reg <= 16'h0C11;
            14'h59 : data_reg <= 16'h211C;
            14'h5A : data_reg <= 16'h1333;
            14'h5B : data_reg <= 16'h0C13;
            14'h5C : data_reg <= 16'hA302;
            14'h5D : data_reg <= 16'h1CE6;
            14'h5E : data_reg <= 16'h1B0D;
            14'h5F : data_reg <= 16'h280C;
            14'h60 : data_reg <= 16'h0D1C;
            14'h61 : data_reg <= 16'h8C9C;
            14'h62 : data_reg <= 16'h1D6D;
            14'h63 : data_reg <= 16'h8C22;
            14'h64 : data_reg <= 16'h1D5D;
            14'h65 : data_reg <= 16'h221D;
            14'h66 : data_reg <= 16'h001C;
            14'h67 : data_reg <= 16'h3C22;
            14'h68 : data_reg <= 16'h1E3E;
            14'h69 : data_reg <= 16'h00AB;
            14'h6A : data_reg <= 16'h3C23;
            14'h6B : data_reg <= 16'h3EE5;
            14'h6C : data_reg <= 16'h1CD0;
            14'h6D : data_reg <= 16'h1D0B;
            14'h6E : data_reg <= 16'hE00C;
            14'h6F : data_reg <= 16'h1CE2;
            14'h70 : data_reg <= 16'h1B0D;
            14'h71 : data_reg <= 16'h280C;
            14'h72 : data_reg <= 16'h0D1C;
            14'h73 : data_reg <= 16'h8C9C;
            14'h74 : data_reg <= 16'h1D6D;
            14'h75 : data_reg <= 16'h8C22;
            14'h76 : data_reg <= 16'h1D5D;
            14'h77 : data_reg <= 16'h221D;
            14'h78 : data_reg <= 16'h001C;
            14'h79 : data_reg <= 16'h3C22;
            14'h7A : data_reg <= 16'h1E3E;
            14'h7B : data_reg <= 16'h0054;
            14'h7C : data_reg <= 16'h3C23;
            14'h7D : data_reg <= 16'h3EE5;
            14'h7E : data_reg <= 16'h1CD0;
            14'h7F : data_reg <= 16'h1D0B;
            14'h80 : data_reg <= 16'hD00C;
            14'h81 : data_reg <= 16'h1C11;
            14'h82 : data_reg <= 16'h1B0D;
            14'h83 : data_reg <= 16'h280C;
            14'h84 : data_reg <= 16'h0D1C;
            14'h85 : data_reg <= 16'h8C9C;
            14'h86 : data_reg <= 16'h1D6D;
            14'h87 : data_reg <= 16'h8C22;
            14'h88 : data_reg <= 16'h1D5D;
            14'h89 : data_reg <= 16'h221D;
            14'h8A : data_reg <= 16'h001C;
            14'h8B : data_reg <= 16'h3C22;
            14'h8C : data_reg <= 16'h1E3E;
            14'h8D : data_reg <= 16'h0056;
            14'h8E : data_reg <= 16'h3C23;
            14'h8F : data_reg <= 16'h3EE5;
            14'h90 : data_reg <= 16'h1CD0;
            14'h91 : data_reg <= 16'h1D0B;
            14'h92 : data_reg <= 16'hD00C;
            14'h93 : data_reg <= 16'h2012;
            14'h94 : data_reg <= 16'hD113;
            14'h95 : data_reg <= 16'h1CE9;
            14'h96 : data_reg <= 16'h3122;
            14'h97 : data_reg <= 16'h0C11;
            14'h98 : data_reg <= 16'h211C;
            14'h99 : data_reg <= 16'h1333;
            14'h9A : data_reg <= 16'h0C13;
            14'h9B : data_reg <= 16'hA302;
            14'h9C : data_reg <= 16'h1CE6;
            14'h9D : data_reg <= 16'h1B0D;
            14'h9E : data_reg <= 16'h280C;
            14'h9F : data_reg <= 16'h0D1C;
            14'hA0 : data_reg <= 16'h8C9C;
            14'hA1 : data_reg <= 16'h1D6D;
            14'hA2 : data_reg <= 16'h8C22;
            14'hA3 : data_reg <= 16'h1D5D;
            14'hA4 : data_reg <= 16'h221D;
            14'hA5 : data_reg <= 16'h001C;
            14'hA6 : data_reg <= 16'h3C22;
            14'hA7 : data_reg <= 16'h1E3E;
            14'hA8 : data_reg <= 16'h0129;
            14'hA9 : data_reg <= 16'h3C23;
            14'hAA : data_reg <= 16'h3EE5;
            14'hAB : data_reg <= 16'h1CD0;
            14'hAC : data_reg <= 16'h1D0B;
            14'hAD : data_reg <= 16'hE00C;
            14'hAE : data_reg <= 16'h1CE2;
            14'hAF : data_reg <= 16'h1B0D;
            14'hB0 : data_reg <= 16'h280C;
            14'hB1 : data_reg <= 16'h0D1C;
            14'hB2 : data_reg <= 16'h8C9C;
            14'hB3 : data_reg <= 16'h1D6D;
            14'hB4 : data_reg <= 16'h8C22;
            14'hB5 : data_reg <= 16'h1D5D;
            14'hB6 : data_reg <= 16'h221D;
            14'hB7 : data_reg <= 16'h001C;
            14'hB8 : data_reg <= 16'h3C22;
            14'hB9 : data_reg <= 16'h1E3E;
            14'hBA : data_reg <= 16'h0054;
            14'hBB : data_reg <= 16'h3C23;
            14'hBC : data_reg <= 16'h3EE5;
            14'hBD : data_reg <= 16'h1CD0;
            14'hBE : data_reg <= 16'h1D0B;
            14'hBF : data_reg <= 16'hD00C;
            14'hC0 : data_reg <= 16'h1C19;
            14'hC1 : data_reg <= 16'h1B0D;
            14'hC2 : data_reg <= 16'h280C;
            14'hC3 : data_reg <= 16'h0D1C;
            14'hC4 : data_reg <= 16'h8C9C;
            14'hC5 : data_reg <= 16'h1D6D;
            14'hC6 : data_reg <= 16'h8C22;
            14'hC7 : data_reg <= 16'h1D5D;
            14'hC8 : data_reg <= 16'h221D;
            14'hC9 : data_reg <= 16'h001C;
            14'hCA : data_reg <= 16'h3C22;
            14'hCB : data_reg <= 16'h1E3E;
            14'hCC : data_reg <= 16'h005A;
            14'hCD : data_reg <= 16'h3C23;
            14'hCE : data_reg <= 16'h3EE5;
            14'hCF : data_reg <= 16'h1CD0;
            14'hD0 : data_reg <= 16'h1D0B;
            14'hD1 : data_reg <= 16'h1A0C;
            14'hD2 : data_reg <= 16'h1126;
            14'hD3 : data_reg <= 16'hE10A;
            14'hD4 : data_reg <= 16'h0D1C;
            14'hD5 : data_reg <= 16'h0C1B;
            14'hD6 : data_reg <= 16'h1C28;
            14'hD7 : data_reg <= 16'h9C0D;
            14'hD8 : data_reg <= 16'h6D8C;
            14'hD9 : data_reg <= 16'h221D;
            14'hDA : data_reg <= 16'h5D8C;
            14'hDB : data_reg <= 16'h1D1D;
            14'hDC : data_reg <= 16'h1C22;
            14'hDD : data_reg <= 16'h3C22;
            14'hDE : data_reg <= 16'h1E3E;
            14'hDF : data_reg <= 16'h0C80;
            14'hE0 : data_reg <= 16'h3C23;
            14'hE1 : data_reg <= 16'h3EE5;
            14'hE2 : data_reg <= 16'h1CD0;
            14'hE3 : data_reg <= 16'h1D0B;
            14'hE4 : data_reg <= 16'h120C;
            14'hE5 : data_reg <= 16'h1102;
            14'hE6 : data_reg <= 16'hE10A;
            14'hE7 : data_reg <= 16'h1C24;
            14'hE8 : data_reg <= 16'h8C20;
            14'hE9 : data_reg <= 16'h2A1C;
            14'hEA : data_reg <= 16'h115C;
            14'hEB : data_reg <= 16'h1C24;
            14'hEC : data_reg <= 16'h8C20;
            14'hED : data_reg <= 16'h2F1C;
            14'hEE : data_reg <= 16'h315C;
            14'hEF : data_reg <= 16'h0A11;
            14'hF0 : data_reg <= 16'h24E1;
            14'hF1 : data_reg <= 16'h261C;
            14'hF2 : data_reg <= 16'h1C8C;
            14'hF3 : data_reg <= 16'h5C24;
            14'hF4 : data_reg <= 16'h2412;
            14'hF5 : data_reg <= 16'h2C1C;
            14'hF6 : data_reg <= 16'h1C8C;
            14'hF7 : data_reg <= 16'h5C28;
            14'hF8 : data_reg <= 16'h32E5;
            14'hF9 : data_reg <= 16'h11E5;
            14'hFA : data_reg <= 16'hE10A;
            14'hFB : data_reg <= 16'h1C24;
            14'hFC : data_reg <= 16'h8C23;
            14'hFD : data_reg <= 16'h221C;
            14'hFE : data_reg <= 16'hE55C;
            14'hFF : data_reg <= 16'hE532;
            14'h100 : data_reg <= 16'h0A11;
            14'h101 : data_reg <= 16'h24E1;
            14'h102 : data_reg <= 16'h2A1C;
            14'h103 : data_reg <= 16'h1C8C;
            14'h104 : data_reg <= 16'h5C2A;
            14'h105 : data_reg <= 16'h2412;
            14'h106 : data_reg <= 16'h251C;
            14'h107 : data_reg <= 16'h1C8C;
            14'h108 : data_reg <= 16'h5C25;
            14'h109 : data_reg <= 16'h1142;
            14'h10A : data_reg <= 16'hE10A;
            14'h10B : data_reg <= 16'h4222;
            14'h10C : data_reg <= 16'h0A11;
            14'h10D : data_reg <= 16'h24E1;
            14'h10E : data_reg <= 16'h2A1C;
            14'h10F : data_reg <= 16'h1C8C;
            14'h110 : data_reg <= 16'h5C2A;
            14'h111 : data_reg <= 16'h2412;
            14'h112 : data_reg <= 16'h251C;
            14'h113 : data_reg <= 16'h1C8C;
            14'h114 : data_reg <= 16'h5C25;
            14'h115 : data_reg <= 16'h1152;
            14'h116 : data_reg <= 16'hE10A;
            14'h117 : data_reg <= 16'h132D;
            14'h118 : data_reg <= 16'h632E;
            14'h119 : data_reg <= 16'h0A11;
            14'h11A : data_reg <= 16'h72E1;
            14'h11B : data_reg <= 16'h0A11;
            14'h11C : data_reg <= 16'h21E1;
            14'h11D : data_reg <= 16'h2712;
            14'h11E : data_reg <= 16'h1182;
            14'h11F : data_reg <= 16'hE10A;
            14'h120 : data_reg <= 16'h9226;
            14'h121 : data_reg <= 16'h0A11;
            14'h122 : data_reg <= 16'h21E1;
            14'h123 : data_reg <= 16'h2111;
            14'h124 : data_reg <= 16'h1CA1;
            14'h125 : data_reg <= 16'h1B0D;
            14'h126 : data_reg <= 16'h280C;
            14'h127 : data_reg <= 16'h0D1C;
            14'h128 : data_reg <= 16'h8C9C;
            14'h129 : data_reg <= 16'h1D6D;
            14'h12A : data_reg <= 16'h8C22;
            14'h12B : data_reg <= 16'h1D5D;
            14'h12C : data_reg <= 16'h221D;
            14'h12D : data_reg <= 16'h001C;
            14'h12E : data_reg <= 16'h3C22;
            14'h12F : data_reg <= 16'h1E3E;
            14'h130 : data_reg <= 16'h028E;
            14'h131 : data_reg <= 16'h3C23;
            14'h132 : data_reg <= 16'h3EE5;
            14'h133 : data_reg <= 16'h1CD0;
            14'h134 : data_reg <= 16'h1D0B;
            14'h135 : data_reg <= 16'hE00C;
            14'h136 : data_reg <= 16'h0D1C;
            14'h137 : data_reg <= 16'h0C1B;
            14'h138 : data_reg <= 16'h1C28;
            14'h139 : data_reg <= 16'h9C0D;
            14'h13A : data_reg <= 16'h6D8C;
            14'h13B : data_reg <= 16'h221D;
            14'h13C : data_reg <= 16'h5D8C;
            14'h13D : data_reg <= 16'h1D1D;
            14'h13E : data_reg <= 16'h1C22;
            14'h13F : data_reg <= 16'h3C22;
            14'h140 : data_reg <= 16'h1E3E;
            14'h141 : data_reg <= 16'h03B8;
            14'h142 : data_reg <= 16'h3C23;
            14'h143 : data_reg <= 16'h3EE5;
            14'h144 : data_reg <= 16'h1CD0;
            14'h145 : data_reg <= 16'h1D0B;
            14'h146 : data_reg <= 16'h1E0C;
            14'h147 : data_reg <= 16'hA120;
            14'h148 : data_reg <= 16'h0D1C;
            14'h149 : data_reg <= 16'h0C1B;
            14'h14A : data_reg <= 16'h1C28;
            14'h14B : data_reg <= 16'h9C0D;
            14'h14C : data_reg <= 16'h6D8C;
            14'h14D : data_reg <= 16'h221D;
            14'h14E : data_reg <= 16'h5D8C;
            14'h14F : data_reg <= 16'h1D1D;
            14'h150 : data_reg <= 16'h1C22;
            14'h151 : data_reg <= 16'h3C22;
            14'h152 : data_reg <= 16'h1E3E;
            14'h153 : data_reg <= 16'h03B8;
            14'h154 : data_reg <= 16'h3C23;
            14'h155 : data_reg <= 16'h3EE5;
            14'h156 : data_reg <= 16'h1CD0;
            14'h157 : data_reg <= 16'h1D0B;
            14'h158 : data_reg <= 16'hE00C;
            14'h159 : data_reg <= 16'hB121;
            14'h15A : data_reg <= 16'h0D1C;
            14'h15B : data_reg <= 16'h0C1B;
            14'h15C : data_reg <= 16'h1C28;
            14'h15D : data_reg <= 16'h9C0D;
            14'h15E : data_reg <= 16'h6D8C;
            14'h15F : data_reg <= 16'h221D;
            14'h160 : data_reg <= 16'h5D8C;
            14'h161 : data_reg <= 16'h1D1D;
            14'h162 : data_reg <= 16'h1C22;
            14'h163 : data_reg <= 16'h3C22;
            14'h164 : data_reg <= 16'h1E3E;
            14'h165 : data_reg <= 16'h03B8;
            14'h166 : data_reg <= 16'h3C23;
            14'h167 : data_reg <= 16'h3EE5;
            14'h168 : data_reg <= 16'h1CD0;
            14'h169 : data_reg <= 16'h1D0B;
            14'h16A : data_reg <= 16'hE00C;
            14'h16B : data_reg <= 16'hB120;
            14'h16C : data_reg <= 16'h0D1C;
            14'h16D : data_reg <= 16'h0C1B;
            14'h16E : data_reg <= 16'h1C28;
            14'h16F : data_reg <= 16'h9C0D;
            14'h170 : data_reg <= 16'h6D8C;
            14'h171 : data_reg <= 16'h221D;
            14'h172 : data_reg <= 16'h5D8C;
            14'h173 : data_reg <= 16'h1D1D;
            14'h174 : data_reg <= 16'h1C22;
            14'h175 : data_reg <= 16'h3C22;
            14'h176 : data_reg <= 16'h1E3E;
            14'h177 : data_reg <= 16'h031C;
            14'h178 : data_reg <= 16'h3C23;
            14'h179 : data_reg <= 16'h3EE5;
            14'h17A : data_reg <= 16'h1CD0;
            14'h17B : data_reg <= 16'h1D0B;
            14'h17C : data_reg <= 16'hE00C;
            14'h17D : data_reg <= 16'h0D1C;
            14'h17E : data_reg <= 16'h0C1B;
            14'h17F : data_reg <= 16'h1C28;
            14'h180 : data_reg <= 16'h9C0D;
            14'h181 : data_reg <= 16'h6D8C;
            14'h182 : data_reg <= 16'h221D;
            14'h183 : data_reg <= 16'h5D8C;
            14'h184 : data_reg <= 16'h1D1D;
            14'h185 : data_reg <= 16'h1C22;
            14'h186 : data_reg <= 16'h3C22;
            14'h187 : data_reg <= 16'h1E3E;
            14'h188 : data_reg <= 16'h03B8;
            14'h189 : data_reg <= 16'h3C23;
            14'h18A : data_reg <= 16'h3EE5;
            14'h18B : data_reg <= 16'h1CD0;
            14'h18C : data_reg <= 16'h1D0B;
            14'h18D : data_reg <= 16'h1E0C;
            14'h18E : data_reg <= 16'h1C24;
            14'h18F : data_reg <= 16'h8C25;
            14'h190 : data_reg <= 16'h2A1C;
            14'h191 : data_reg <= 16'hCF5C;
            14'h192 : data_reg <= 16'hDF20;
            14'h193 : data_reg <= 16'h0A11;
            14'h194 : data_reg <= 16'h24E1;
            14'h195 : data_reg <= 16'h251C;
            14'h196 : data_reg <= 16'h1C8C;
            14'h197 : data_reg <= 16'h5C20;
            14'h198 : data_reg <= 16'h20E4;
            14'h199 : data_reg <= 16'h11E3;
            14'h19A : data_reg <= 16'hE10A;
            14'h19B : data_reg <= 16'h1C24;
            14'h19C : data_reg <= 16'h8C20;
            14'h19D : data_reg <= 16'h2D1C;
            14'h19E : data_reg <= 16'hE55C;
            14'h19F : data_reg <= 16'h0A11;
            14'h1A0 : data_reg <= 16'h1CE1;
            14'h1A1 : data_reg <= 16'h1B0D;
            14'h1A2 : data_reg <= 16'h280C;
            14'h1A3 : data_reg <= 16'h0D1C;
            14'h1A4 : data_reg <= 16'h8C9C;
            14'h1A5 : data_reg <= 16'h1D6D;
            14'h1A6 : data_reg <= 16'h8C22;
            14'h1A7 : data_reg <= 16'h1D5D;
            14'h1A8 : data_reg <= 16'h221D;
            14'h1A9 : data_reg <= 16'h001C;
            14'h1AA : data_reg <= 16'h3C22;
            14'h1AB : data_reg <= 16'h1E3E;
            14'h1AC : data_reg <= 16'h03B9;
            14'h1AD : data_reg <= 16'h3C23;
            14'h1AE : data_reg <= 16'h3EE5;
            14'h1AF : data_reg <= 16'h1CD0;
            14'h1B0 : data_reg <= 16'h1D0B;
            14'h1B1 : data_reg <= 16'hE10C;
            14'h1B2 : data_reg <= 16'h1121;
            14'h1B3 : data_reg <= 16'hA121;
            14'h1B4 : data_reg <= 16'h0D1C;
            14'h1B5 : data_reg <= 16'h0C1B;
            14'h1B6 : data_reg <= 16'h1C28;
            14'h1B7 : data_reg <= 16'h9C0D;
            14'h1B8 : data_reg <= 16'h6D8C;
            14'h1B9 : data_reg <= 16'h221D;
            14'h1BA : data_reg <= 16'h5D8C;
            14'h1BB : data_reg <= 16'h1D1D;
            14'h1BC : data_reg <= 16'h1C22;
            14'h1BD : data_reg <= 16'h3C22;
            14'h1BE : data_reg <= 16'h1E3E;
            14'h1BF : data_reg <= 16'h03B8;
            14'h1C0 : data_reg <= 16'h3C23;
            14'h1C1 : data_reg <= 16'h3EE5;
            14'h1C2 : data_reg <= 16'h1CD0;
            14'h1C3 : data_reg <= 16'h1D0B;
            14'h1C4 : data_reg <= 16'hE60C;
            14'h1C5 : data_reg <= 16'h28E0;
            14'h1C6 : data_reg <= 16'h113F;
            14'h1C7 : data_reg <= 16'h0D1C;
            14'h1C8 : data_reg <= 16'h0C1B;
            14'h1C9 : data_reg <= 16'h1C28;
            14'h1CA : data_reg <= 16'h9C0D;
            14'h1CB : data_reg <= 16'h6D8C;
            14'h1CC : data_reg <= 16'h221D;
            14'h1CD : data_reg <= 16'h5D8C;
            14'h1CE : data_reg <= 16'h1D1D;
            14'h1CF : data_reg <= 16'h1C22;
            14'h1D0 : data_reg <= 16'h3C22;
            14'h1D1 : data_reg <= 16'h1E3E;
            14'h1D2 : data_reg <= 16'hFFFF;
            14'h1D3 : data_reg <= 16'h3C23;
            14'h1D4 : data_reg <= 16'h3EE5;
            14'h1D5 : data_reg <= 16'h1CD0;
            14'h1D6 : data_reg <= 16'h1D0B;
            14'h1D7 : data_reg <= 16'hE70C;
            14'h1D8 : data_reg <= 16'h20C1;
            14'h1D9 : data_reg <= 16'hE7D1;
            14'h1DA : data_reg <= 16'h0A11;
            14'h1DB : data_reg <= 16'hE2E1;
            14'h1DC : data_reg <= 16'h2AE8;
            14'h1DD : data_reg <= 16'h0A11;
            14'h1DE : data_reg <= 16'hE2E1;
            14'h1DF : data_reg <= 16'h0D1C;
            14'h1E0 : data_reg <= 16'h0C1B;
            14'h1E1 : data_reg <= 16'h1C28;
            14'h1E2 : data_reg <= 16'h9C0D;
            14'h1E3 : data_reg <= 16'h6D8C;
            14'h1E4 : data_reg <= 16'h221D;
            14'h1E5 : data_reg <= 16'h5D8C;
            14'h1E6 : data_reg <= 16'h1D1D;
            14'h1E7 : data_reg <= 16'h1C22;
            14'h1E8 : data_reg <= 16'h3C22;
            14'h1E9 : data_reg <= 16'h1E3E;
            14'h1EA : data_reg <= 16'h0058;
            14'h1EB : data_reg <= 16'h3C23;
            14'h1EC : data_reg <= 16'h3EE5;
            14'h1ED : data_reg <= 16'h1CD0;
            14'h1EE : data_reg <= 16'h1D0B;
            14'h1EF : data_reg <= 16'hD00C;
            14'h1F0 : data_reg <= 16'h1C1F;
            14'h1F1 : data_reg <= 16'h1B0D;
            14'h1F2 : data_reg <= 16'h280C;
            14'h1F3 : data_reg <= 16'h0D1C;
            14'h1F4 : data_reg <= 16'h8C9C;
            14'h1F5 : data_reg <= 16'h1D6D;
            14'h1F6 : data_reg <= 16'h8C22;
            14'h1F7 : data_reg <= 16'h1D5D;
            14'h1F8 : data_reg <= 16'h221D;
            14'h1F9 : data_reg <= 16'h001C;
            14'h1FA : data_reg <= 16'h3C22;
            14'h1FB : data_reg <= 16'h1E3E;
            14'h1FC : data_reg <= 16'h0062;
            14'h1FD : data_reg <= 16'h3C23;
            14'h1FE : data_reg <= 16'h3EE5;
            14'h1FF : data_reg <= 16'h1CD0;
            14'h200 : data_reg <= 16'h1D0B;
            14'h201 : data_reg <= 16'hE10C;
            14'h202 : data_reg <= 16'h0D1C;
            14'h203 : data_reg <= 16'h0C1B;
            14'h204 : data_reg <= 16'h1C28;
            14'h205 : data_reg <= 16'h9C0D;
            14'h206 : data_reg <= 16'h6D8C;
            14'h207 : data_reg <= 16'h221D;
            14'h208 : data_reg <= 16'h5D8C;
            14'h209 : data_reg <= 16'h1D1D;
            14'h20A : data_reg <= 16'h1C22;
            14'h20B : data_reg <= 16'h3C22;
            14'h20C : data_reg <= 16'h1E3E;
            14'h20D : data_reg <= 16'h015D;
            14'h20E : data_reg <= 16'h3C23;
            14'h20F : data_reg <= 16'h3EE5;
            14'h210 : data_reg <= 16'h1CD0;
            14'h211 : data_reg <= 16'h1D0B;
            14'h212 : data_reg <= 16'hE10C;
            14'h213 : data_reg <= 16'h0D1C;
            14'h214 : data_reg <= 16'h0C1B;
            14'h215 : data_reg <= 16'h1C28;
            14'h216 : data_reg <= 16'h9C0D;
            14'h217 : data_reg <= 16'h6D8C;
            14'h218 : data_reg <= 16'h221D;
            14'h219 : data_reg <= 16'h5D8C;
            14'h21A : data_reg <= 16'h1D1D;
            14'h21B : data_reg <= 16'h1C22;
            14'h21C : data_reg <= 16'h3C22;
            14'h21D : data_reg <= 16'h1E3E;
            14'h21E : data_reg <= 16'h00DF;
            14'h21F : data_reg <= 16'h3C23;
            14'h220 : data_reg <= 16'h3EE5;
            14'h221 : data_reg <= 16'h1CD0;
            14'h222 : data_reg <= 16'h1D0B;
            14'h223 : data_reg <= 16'hE10C;
            14'h224 : data_reg <= 16'h00E8;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
