module rom05(input clk, input enable, input [30-1:0] addr, output [32-1:0] data);
    reg [32-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            30'h0 : data_reg <= 32'h4D525341;
            30'h1 : data_reg <= 32'h9C0D1C28;
            30'h2 : data_reg <= 32'h231D6D8C;
            30'h3 : data_reg <= 32'h1C1D5D8C;
            30'h4 : data_reg <= 32'h280C1B0D;
            30'h5 : data_reg <= 32'h8C9C0D1C;
            30'h6 : data_reg <= 32'h8C231D6D;
            30'h7 : data_reg <= 32'h241D1D5D;
            30'h8 : data_reg <= 32'h0000001C;
            30'h9 : data_reg <= 32'h1E3E3C22;
            30'hA : data_reg <= 32'h00001000;
            30'hB : data_reg <= 32'h3EE53C23;
            30'hC : data_reg <= 32'h1D0B1CD0;
            30'hD : data_reg <= 32'h0D1C110C;
            30'hE : data_reg <= 32'h1C280C1B;
            30'hF : data_reg <= 32'h6D8C9C0D;
            30'h10 : data_reg <= 32'h5D8C231D;
            30'h11 : data_reg <= 32'h1C241D1D;
            30'h12 : data_reg <= 32'h1E3E3C22;
            30'h13 : data_reg <= 32'hABCDEF00;
            30'h14 : data_reg <= 32'h3EE53C23;
            30'h15 : data_reg <= 32'h1D0B1CD0;
            30'h16 : data_reg <= 32'h0D1C120C;
            30'h17 : data_reg <= 32'h1C280C1B;
            30'h18 : data_reg <= 32'h6D8C9C0D;
            30'h19 : data_reg <= 32'h5D8C231D;
            30'h1A : data_reg <= 32'h1C241D1D;
            30'h1B : data_reg <= 32'h1E3E3C22;
            30'h1C : data_reg <= 32'h01020304;
            30'h1D : data_reg <= 32'h3EE53C23;
            30'h1E : data_reg <= 32'h1D0B1CD0;
            30'h1F : data_reg <= 32'h0D1C130C;
            30'h20 : data_reg <= 32'h1C280C1B;
            30'h21 : data_reg <= 32'h6D8C9C0D;
            30'h22 : data_reg <= 32'h5D8C231D;
            30'h23 : data_reg <= 32'h1C241D1D;
            30'h24 : data_reg <= 32'h1E3E3C22;
            30'h25 : data_reg <= 32'h0000012B;
            30'h26 : data_reg <= 32'h3EE53C23;
            30'h27 : data_reg <= 32'h1D0B1CD0;
            30'h28 : data_reg <= 32'h1C24EC0C;
            30'h29 : data_reg <= 32'h221C8C22;
            30'h2A : data_reg <= 32'hC1021D5C;
            30'h2B : data_reg <= 32'h03113124;
            30'h2C : data_reg <= 32'h113124C1;
            30'h2D : data_reg <= 32'h9C0D1C28;
            30'h2E : data_reg <= 32'h221D6D8C;
            30'h2F : data_reg <= 32'h021D5D8C;
            30'h30 : data_reg <= 32'h113122C1;
            30'h31 : data_reg <= 32'h3122C103;
            30'h32 : data_reg <= 32'h0D1C2811;
            30'h33 : data_reg <= 32'h1D6D8C9C;
            30'h34 : data_reg <= 32'h1D5D8C21;
            30'h35 : data_reg <= 32'h3121C12A;
            30'h36 : data_reg <= 32'h21C12B11;
            30'h37 : data_reg <= 32'hC12C1131;
            30'h38 : data_reg <= 32'h2D113121;
            30'h39 : data_reg <= 32'h113121C1;
            30'h3A : data_reg <= 32'h9C0D1C28;
            30'h3B : data_reg <= 32'h231D6D8C;
            30'h3C : data_reg <= 32'h1C1D5D8C;
            30'h3D : data_reg <= 32'h280C1B0D;
            30'h3E : data_reg <= 32'h8C9C0D1C;
            30'h3F : data_reg <= 32'h8C231D6D;
            30'h40 : data_reg <= 32'h241D1D5D;
            30'h41 : data_reg <= 32'h0000001C;
            30'h42 : data_reg <= 32'h1E3E3C22;
            30'h43 : data_reg <= 32'h00001000;
            30'h44 : data_reg <= 32'h3EE53C23;
            30'h45 : data_reg <= 32'h1D0B1CD0;
            30'h46 : data_reg <= 32'hE9D1110C;
            30'h47 : data_reg <= 32'hD1113124;
            30'h48 : data_reg <= 32'h113124E9;
            30'h49 : data_reg <= 32'h3124E9D1;
            30'h4A : data_reg <= 32'hE8E9D111;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
