module rom08(input clk, input enable, input [15-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            15'h0 : data_reg <= 16'h5341;
            15'h1 : data_reg <= 16'h4D52;
            15'h2 : data_reg <= 16'h1C28;
            15'h3 : data_reg <= 16'h9C0D;
            15'h4 : data_reg <= 16'h6D8C;
            15'h5 : data_reg <= 16'h211D;
            15'h6 : data_reg <= 16'h5D8C;
            15'h7 : data_reg <= 16'h0D1D;
            15'h8 : data_reg <= 16'h281B;
            15'h9 : data_reg <= 16'h0D1C;
            15'hA : data_reg <= 16'h8C9C;
            15'hB : data_reg <= 16'h1D6D;
            15'hC : data_reg <= 16'h8C21;
            15'hD : data_reg <= 16'h1D5D;
            15'hE : data_reg <= 16'h1C21;
            15'hF : data_reg <= 16'h3C22;
            15'h10 : data_reg <= 16'h1E3E;
            15'h11 : data_reg <= 16'h2355;
            15'h12 : data_reg <= 16'hE53C;
            15'h13 : data_reg <= 16'hD03E;
            15'h14 : data_reg <= 16'h0B1C;
            15'h15 : data_reg <= 16'h0C1D;
            15'h16 : data_reg <= 16'hFD1E;
            15'h17 : data_reg <= 16'h1C24;
            15'h18 : data_reg <= 16'h8C2A;
            15'h19 : data_reg <= 16'h2A1C;
            15'h1A : data_reg <= 16'hEB5C;
            15'h1B : data_reg <= 16'h1B0D;
            15'h1C : data_reg <= 16'h1C28;
            15'h1D : data_reg <= 16'h9C0D;
            15'h1E : data_reg <= 16'h6D8C;
            15'h1F : data_reg <= 16'h211D;
            15'h20 : data_reg <= 16'h5D8C;
            15'h21 : data_reg <= 16'h211D;
            15'h22 : data_reg <= 16'h221C;
            15'h23 : data_reg <= 16'h3E3C;
            15'h24 : data_reg <= 16'h951E;
            15'h25 : data_reg <= 16'h3C23;
            15'h26 : data_reg <= 16'h3EE5;
            15'h27 : data_reg <= 16'h1CD0;
            15'h28 : data_reg <= 16'h1D0B;
            15'h29 : data_reg <= 16'hFA0C;
            15'h2A : data_reg <= 16'h0DEB;
            15'h2B : data_reg <= 16'h281B;
            15'h2C : data_reg <= 16'h0D1C;
            15'h2D : data_reg <= 16'h8C9C;
            15'h2E : data_reg <= 16'h1D6D;
            15'h2F : data_reg <= 16'h8C21;
            15'h30 : data_reg <= 16'h1D5D;
            15'h31 : data_reg <= 16'h1C21;
            15'h32 : data_reg <= 16'h3C22;
            15'h33 : data_reg <= 16'h1E3E;
            15'h34 : data_reg <= 16'h232D;
            15'h35 : data_reg <= 16'hE53C;
            15'h36 : data_reg <= 16'hD03E;
            15'h37 : data_reg <= 16'h0B1C;
            15'h38 : data_reg <= 16'h0C1D;
            15'h39 : data_reg <= 16'h0DEE;
            15'h3A : data_reg <= 16'h281B;
            15'h3B : data_reg <= 16'h0D1C;
            15'h3C : data_reg <= 16'h8C9C;
            15'h3D : data_reg <= 16'h1D6D;
            15'h3E : data_reg <= 16'h8C21;
            15'h3F : data_reg <= 16'h1D5D;
            15'h40 : data_reg <= 16'h1C21;
            15'h41 : data_reg <= 16'h3C22;
            15'h42 : data_reg <= 16'h1E3E;
            15'h43 : data_reg <= 16'h2336;
            15'h44 : data_reg <= 16'hE53C;
            15'h45 : data_reg <= 16'hD03E;
            15'h46 : data_reg <= 16'h0B1C;
            15'h47 : data_reg <= 16'h0C1D;
            15'h48 : data_reg <= 16'h2CED;
            15'h49 : data_reg <= 16'hFE1D;
            15'h4A : data_reg <= 16'hE9E8;
            15'h4B : data_reg <= 16'h00E8;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
