../reflet.vh